
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_mux21_nbit is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_mux21_nbit;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_15 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_15;

architecture SYN_df_nand of mux21_15 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_14 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_14;

architecture SYN_df_nand of mux21_14 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_13 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_13;

architecture SYN_df_nand of mux21_13 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_12 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_12;

architecture SYN_df_nand of mux21_12 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_11 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_11;

architecture SYN_df_nand of mux21_11 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_10 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_10;

architecture SYN_df_nand of mux21_10 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_9 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_9;

architecture SYN_df_nand of mux21_9 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_8 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_8;

architecture SYN_df_nand of mux21_8 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_7 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_7;

architecture SYN_df_nand of mux21_7 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_6 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_6;

architecture SYN_df_nand of mux21_6 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_5 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_5;

architecture SYN_df_nand of mux21_5 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_4 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_4;

architecture SYN_df_nand of mux21_4 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_3 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_3;

architecture SYN_df_nand of mux21_3 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_2 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_2;

architecture SYN_df_nand of mux21_2 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_1 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_1;

architecture SYN_df_nand of mux21_1 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_0 is

   port( x, y, s : in std_logic;  m : out std_logic);

end mux21_0;

architecture SYN_df_nand of mux21_0 is

   component SAEDRVT14_MUX2_MM_0P5
      port( D0, D1, S : in std_logic;  X : out std_logic);
   end component;

begin
   
   U1 : SAEDRVT14_MUX2_MM_0P5 port map( D0 => x, D1 => y, S => s, X => m);

end SYN_df_nand;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_nbit.all;

entity mux21_nbit is

   port( X, y : in std_logic_vector (15 downto 0);  s : in std_logic;  m : out 
         std_logic_vector (15 downto 0));

end mux21_nbit;

architecture SYN_df of mux21_nbit is

   component mux21_1
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_2
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_3
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_4
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_5
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_6
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_7
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_8
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_9
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_10
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_11
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_12
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_13
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_14
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_15
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;
   
   component mux21_0
      port( x, y, s : in std_logic;  m : out std_logic);
   end component;

begin
   
   mux21_i_0 : mux21_0 port map( x => X(0), y => y(0), s => s, m => m(0));
   mux21_i_1 : mux21_15 port map( x => X(1), y => y(1), s => s, m => m(1));
   mux21_i_2 : mux21_14 port map( x => X(2), y => y(2), s => s, m => m(2));
   mux21_i_3 : mux21_13 port map( x => X(3), y => y(3), s => s, m => m(3));
   mux21_i_4 : mux21_12 port map( x => X(4), y => y(4), s => s, m => m(4));
   mux21_i_5 : mux21_11 port map( x => X(5), y => y(5), s => s, m => m(5));
   mux21_i_6 : mux21_10 port map( x => X(6), y => y(6), s => s, m => m(6));
   mux21_i_7 : mux21_9 port map( x => X(7), y => y(7), s => s, m => m(7));
   mux21_i_8 : mux21_8 port map( x => X(8), y => y(8), s => s, m => m(8));
   mux21_i_9 : mux21_7 port map( x => X(9), y => y(9), s => s, m => m(9));
   mux21_i_10 : mux21_6 port map( x => X(10), y => y(10), s => s, m => m(10));
   mux21_i_11 : mux21_5 port map( x => X(11), y => y(11), s => s, m => m(11));
   mux21_i_12 : mux21_4 port map( x => X(12), y => y(12), s => s, m => m(12));
   mux21_i_13 : mux21_3 port map( x => X(13), y => y(13), s => s, m => m(13));
   mux21_i_14 : mux21_2 port map( x => X(14), y => y(14), s => s, m => m(14));
   mux21_i_15 : mux21_1 port map( x => X(15), y => y(15), s => s, m => m(15));

end SYN_df;
