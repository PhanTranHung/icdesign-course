** Voltage divider **

R1 in out 1K
R2 out 0 1K
V1 in 0  DC 4V
.OP
.END